import EPI_pkg::*;

module segre_tlb (
    input clk_i,
    input rsn_i
);


endmodule : segre_tlb
